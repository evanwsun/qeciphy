// SPDX-License-Identifier: LicenseRef-LICENSE
// -----------------------------------------------------------------------------
// File        : qeciphy_clk_mmcm.sv
// Description : Lint stub for Xilinx clocking wizard module.
//               Declares the module interface for tooling convenience only.
//               No functional implementation is provided.
// 
// Copyright (c) 2025 Riverlane Ltd.
// This file is not affiliated with or endorsed by Xilinx Inc. or AMD.
// The module names and ports are reproduced solely for build compatibility.
// -----------------------------------------------------------------------------

module qeciphy_clk_mmcm (
    output clk_out_2x,
    output clk_out,
    input  reset,
    output input_clk_stopped,
    input  clk_in
);

endmodule
